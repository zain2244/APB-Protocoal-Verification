///`include "interface.sv"
`include "transaction.sv"
`include "apb_config.sv"
`include "seq_case.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "enviroment.sv"